-- 32 = ' '
32*8+0 => b"00000000"
32*8+1 => b"00000000"
32*8+2 => b"00000000"
32*8+3 => b"00000000"
32*8+4 => b"00000000"
32*8+5 => b"00000000"
32*8+6 => b"00000000"
32*8+7 => b"00000000"

-- 37 = '%'
37*8+0 => b"00000000"
37*8+1 => b"00100010"
37*8+2 => b"01010100"
37*8+3 => b"00101000"
37*8+4 => b"00001010"
37*8+5 => b"00010101"
37*8+6 => b"00100010"
37*8+7 => b"00000000"

-- 42 = '*'
42*8+0 => b"00000000"
42*8+1 => b"00000000"
42*8+2 => b"00010000"
42*8+3 => b"01010100"
42*8+4 => b"00101000"
42*8+5 => b"01010100"
42*8+6 => b"00010000"
42*8+7 => b"00000000"

-- 43 = '+'
43*8+0 => b"00000000"
43*8+1 => b"00010000"
43*8+2 => b"00010000"
43*8+3 => b"01111100"
43*8+4 => b"00010000"
43*8+5 => b"00010000"
43*8+6 => b"00000000"
43*8+7 => b"00000000"

-- 45 = '-'
45*8+0 => b"00000000"
45*8+1 => b"00000000"
45*8+2 => b"00000000"
45*8+3 => b"01111100"
45*8+4 => b"00000000"
45*8+5 => b"00000000"
45*8+6 => b"00000000"
45*8+7 => b"00000000"

-- 46 = '.'
46*8+0 => b"00000000"
46*8+1 => b"00011000"
46*8+2 => b"00111100"
46*8+3 => b"01111110"
46*8+4 => b"01111110"
46*8+5 => b"00111100"
46*8+6 => b"00011000"
46*8+7 => b"00000000"

-- 47 = '/'
47*8+0 => b"00000000"
47*8+1 => b"00000100"
47*8+2 => b"00001000"
47*8+3 => b"00010000"
47*8+4 => b"00100000"
47*8+5 => b"01000000"
47*8+6 => b"00000000"
47*8+7 => b"00000000"

-- 48 = '0'
48*8+0 => b"00111100"
48*8+1 => b"01000110"
48*8+2 => b"01001010"
48*8+3 => b"01001010"
48*8+4 => b"01010010"
48*8+5 => b"01100010"
48*8+6 => b"00111100"
48*8+7 => b"00000000"

-- 49 = '1'
49*8+0 => b"00010000"
49*8+1 => b"00110000"
49*8+2 => b"01110000"
49*8+3 => b"00010000"
49*8+4 => b"00010000"
49*8+5 => b"00010000"
49*8+6 => b"01111100"
49*8+7 => b"00000000"

-- 50 = '2'
50*8+0 => b"00111000"
50*8+1 => b"01000100"
50*8+2 => b"00000100"
50*8+3 => b"00001000"
50*8+4 => b"00010000"
50*8+5 => b"00100000"
50*8+6 => b"01111100"
50*8+7 => b"00000000"

-- 51 = '3'
51*8+0 => b"00111000"
51*8+1 => b"01000100"
51*8+2 => b"00000100"
51*8+3 => b"00111000"
51*8+4 => b"00000100"
51*8+5 => b"01000100"
51*8+6 => b"00111000"
51*8+7 => b"00000000"

-- 52 = '4'
52*8+0 => b"01000100"
52*8+1 => b"01000100"
52*8+2 => b"01000100"
52*8+3 => b"01111100"
52*8+4 => b"00000100"
52*8+5 => b"00000100"
52*8+6 => b"00000100"
52*8+7 => b"00000000"

-- 53 = '5'
53*8+0 => b"01111100"
53*8+1 => b"01000000"
53*8+2 => b"01000000"
53*8+3 => b"01111000"
53*8+4 => b"00000100"
53*8+5 => b"00000100"
53*8+6 => b"01111100"
53*8+7 => b"00000000"

-- 54 = '6'
54*8+0 => b"00111100"
54*8+1 => b"01000000"
54*8+2 => b"01000000"
54*8+3 => b"01111100"
54*8+4 => b"01000010"
54*8+5 => b"01000010"
54*8+6 => b"00111100"
54*8+7 => b"00000000"

-- 55 = '7'
55*8+0 => b"01111110"
55*8+1 => b"00000010"
55*8+2 => b"00000100"
55*8+3 => b"00011100"
55*8+4 => b"00010000"
55*8+5 => b"00100000"
55*8+6 => b"01000000"
55*8+7 => b"00000000"

-- 56 = '8'
56*8+0 => b"00111100"
56*8+1 => b"01000010"
56*8+2 => b"01000010"
56*8+3 => b"00111100"
56*8+4 => b"01000010"
56*8+5 => b"01000010"
56*8+6 => b"00111100"
56*8+7 => b"00000000"

-- 57 = '9'
57*8+0 => b"00111100"
57*8+1 => b"01000010"
57*8+2 => b"01000010"
57*8+3 => b"00111110"
57*8+4 => b"00000010"
57*8+5 => b"00000010"
57*8+6 => b"01111100"
57*8+7 => b"00000000"

-- 60 = '<'
60*8+0 => b"00000000"
60*8+1 => b"00001100"
60*8+2 => b"00010000"
60*8+3 => b"00100000"
60*8+4 => b"00010000"
60*8+5 => b"00001100"
60*8+6 => b"00000000"
60*8+7 => b"00000000"

-- 61 = '='
61*8+0 => b"00000000"
61*8+1 => b"00000000"
61*8+2 => b"01111100"
61*8+3 => b"00000000"
61*8+4 => b"00000000"
61*8+5 => b"01111100"
61*8+6 => b"00000000"
61*8+7 => b"00000000"

-- 62 = '>'
62*8+0 => b"00000000"
62*8+1 => b"00110000"
62*8+2 => b"00001000"
62*8+3 => b"00000100"
62*8+4 => b"00001000"
62*8+5 => b"00110000"
62*8+6 => b"00000000"
62*8+7 => b"00000000"

-- 65 = 'A'
65*8+0 => b"00111000"
65*8+1 => b"01000100"
65*8+2 => b"01000100"
65*8+3 => b"01000100"
65*8+4 => b"01111100"
65*8+5 => b"01000100"
65*8+6 => b"01000100"
65*8+7 => b"00000000"

-- 66 = 'B'
66*8+0 => b"01111000"
66*8+1 => b"01000100"
66*8+2 => b"01000100"
66*8+3 => b"01111000"
66*8+4 => b"01000100"
66*8+5 => b"01000100"
66*8+6 => b"01111000"
66*8+7 => b"00000000"

-- 67 = 'C'
67*8+0 => b"00011100"
67*8+1 => b"00100000"
67*8+2 => b"01000000"
67*8+3 => b"01000000"
67*8+4 => b"01000000"
67*8+5 => b"00100000"
67*8+6 => b"00011100"
67*8+7 => b"00000000"

-- 68 = 'D'
68*8+0 => b"01111000"
68*8+1 => b"01000100"
68*8+2 => b"01000010"
68*8+3 => b"01000010"
68*8+4 => b"01000010"
68*8+5 => b"01000100"
68*8+6 => b"01111000"
68*8+7 => b"00000000"

-- 69 = 'E'
69*8+0 => b"01111100"
69*8+1 => b"01000000"
69*8+2 => b"01000000"
69*8+3 => b"01111100"
69*8+4 => b"01000000"
69*8+5 => b"01000000"
69*8+6 => b"01111100"
69*8+7 => b"00000000"

-- 70 = 'F'
70*8+0 => b"01111100"
70*8+1 => b"01000000"
70*8+2 => b"01000000"
70*8+3 => b"01111100"
70*8+4 => b"01000000"
70*8+5 => b"01000000"
70*8+6 => b"01000000"
70*8+7 => b"00000000"

-- 71 = 'G'
71*8+0 => b"00011100"
71*8+1 => b"00100010"
71*8+2 => b"01000000"
71*8+3 => b"01000110"
71*8+4 => b"01000010"
71*8+5 => b"00100010"
71*8+6 => b"00011100"
71*8+7 => b"00000000"

-- 72 = 'H'
72*8+0 => b"01000010"
72*8+1 => b"01000010"
72*8+2 => b"01000010"
72*8+3 => b"01111110"
72*8+4 => b"01000010"
72*8+5 => b"01000010"
72*8+6 => b"01000010"
72*8+7 => b"00000000"

-- 73 = 'I'
73*8+0 => b"00111000"
73*8+1 => b"00010000"
73*8+2 => b"00010000"
73*8+3 => b"00010000"
73*8+4 => b"00010000"
73*8+5 => b"00010000"
73*8+6 => b"00111000"
73*8+7 => b"00000000"

-- 74 = 'J'
74*8+0 => b"01111110"
74*8+1 => b"00001000"
74*8+2 => b"00001000"
74*8+3 => b"00001000"
74*8+4 => b"00001000"
74*8+5 => b"00001000"
74*8+6 => b"00110000"
74*8+7 => b"00000000"

-- 75 = 'K'
75*8+0 => b"01000000"
75*8+1 => b"01001100"
75*8+2 => b"01010000"
75*8+3 => b"01100000"
75*8+4 => b"01010000"
75*8+5 => b"01001000"
75*8+6 => b"01000100"
75*8+7 => b"00000000"

-- 76 = 'L'
76*8+0 => b"01000000"
76*8+1 => b"01000000"
76*8+2 => b"01000000"
76*8+3 => b"01000000"
76*8+4 => b"01000000"
76*8+5 => b"01000000"
76*8+6 => b"01111000"
76*8+7 => b"00000000"

-- 78 = 'N'
78*8+0 => b"01000010"
78*8+1 => b"01100010"
78*8+2 => b"01010010"
78*8+3 => b"01010010"
78*8+4 => b"01001010"
78*8+5 => b"01000110"
78*8+6 => b"01000010"
78*8+7 => b"00000000"

-- 79 = 'O'
79*8+0 => b"00111000"
79*8+1 => b"01000100"
79*8+2 => b"01000100"
79*8+3 => b"01000100"
79*8+4 => b"01000100"
79*8+5 => b"01000100"
79*8+6 => b"00111000"
79*8+7 => b"00000000"

-- 80 = 'P'
80*8+0 => b"01111000"
80*8+1 => b"01000100"
80*8+2 => b"01000100"
80*8+3 => b"01111000"
80*8+4 => b"01000000"
80*8+5 => b"01000000"
80*8+6 => b"01000000"
80*8+7 => b"00000000"

-- 82 = 'R'
82*8+0 => b"01111000"
82*8+1 => b"01000100"
82*8+2 => b"01000100"
82*8+3 => b"01111000"
82*8+4 => b"01001000"
82*8+5 => b"01001000"
82*8+6 => b"01000100"
82*8+7 => b"00000000"

-- 83 = 'S'
83*8+0 => b"00111000"
83*8+1 => b"01000000"
83*8+2 => b"01000000"
83*8+3 => b"00111000"
83*8+4 => b"00000100"
83*8+5 => b"00000100"
83*8+6 => b"00111000"
83*8+7 => b"00000000"

-- 84 = 'T'
84*8+0 => b"01111100"
84*8+1 => b"00010000"
84*8+2 => b"00010000"
84*8+3 => b"00010000"
84*8+4 => b"00010000"
84*8+5 => b"00010000"
84*8+6 => b"00010000"
84*8+7 => b"00000000"

-- 85 = 'U'
85*8+0 => b"01000010"
85*8+1 => b"01000010"
85*8+2 => b"01000010"
85*8+3 => b"01000010"
85*8+4 => b"01000010"
85*8+5 => b"01000010"
85*8+6 => b"00111100"
85*8+7 => b"00000000"

-- 86 = 'V'
86*8+0 => b"01000010"
86*8+1 => b"01000010"
86*8+2 => b"01000010"
86*8+3 => b"01000010"
86*8+4 => b"01000010"
86*8+5 => b"00100100"
86*8+6 => b"00011000"
86*8+7 => b"00000000"

-- 88 = 'X'
88*8+0 => b"01000100"
88*8+1 => b"01000100"
88*8+2 => b"00101000"
88*8+3 => b"00010000"
88*8+4 => b"00101000"
88*8+6 => b"01000100"
88*8+7 => b"00000000"

-- 89 = 'Y'
89*8+0 => b"01000100"
89*8+1 => b"01000100"
89*8+2 => b"01000100"
89*8+3 => b"00111000"
89*8+4 => b"00010000"
89*8+5 => b"00010000"
89*8+6 => b"00010000"
89*8+7 => b"00000000"

-- 95 = '_'
95*8+0 => b"00000000"
95*8+1 => b"00000000"
95*8+2 => b"00000000"
95*8+3 => b"00000000"
95*8+4 => b"00000000"
95*8+5 => b"00000000"
95*8+6 => b"01111100"
95*8+7 => b"00000000"

-- 120 = BLOCK
120*8+0 => b"11111111"
120*8+1 => b"11111111"
120*8+2 => b"11111111"
120*8+3 => b"11111111"
120*8+4 => b"11111111"
120*8+5 => b"11111111"
120*8+6 => b"11111111"
120*8+7 => b"11111111"
